module B16X4 (
    input wire [15:0] a,
    output wire [3:0] AN,
    output wire [63:0] DISPLAY);



endmodule

// module OneTwoDec (
//     input s,
//     output [1:0] o
// );
//     o[0] = 0;
//     s == 1 ? o[1] = 1 : o[1] = 0;
// endmodule
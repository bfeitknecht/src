module FourOneMux(

);
    
endmodule
module FullAdder (input a, input b, input ci, output s, output co);

endmodule
module Top(
    input [1:0] s,
    output [3:0] AN
);

endmodule
```
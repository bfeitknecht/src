module TwoFourDec (
    input [1:0] s,
    output [3:0] o
);
    
    
endmodule
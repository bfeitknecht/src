module FORD(

);

endmodule
module TwoOneMux(
    input a,
    input b,
    input sel,
    output o
);

endmodule
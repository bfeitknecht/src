module Arithmetic (

)
endmodule
module hw;
  initial
    begin
      $display("Hello, World");
      $finish ;
    end
endmodule
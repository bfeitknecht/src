module FSM (
    input clk,
    input reset,
    input enable,
    output A, B, C
    );

    reg [2:0] state_prev, state_next;

    parameter S0 = 3'b000;
    parameter S1 = 3'b001;
    parameter S2 = 3'b011;
    parameter S3 = 3'b111;

    // state holding register
    always @ (posedge clk, posedge reset) begin
        if (reset == '1') state_prev <= S0;
        else state_prev <= state_next;
    end

    // next state logic 
    always @ (*) begin
        case (state_prev)
            S0: state_next <= (enable == '1') ? S1 : S0;
            S1: state_next <= S2;
            S2: state_next <= S3;
            S3: state_next <= S0;
        endcase
    end

    // output logic
    assign {A, B, C} = state_prev;
endmodule


/*
S0
S1
S2
S3
*/
module Logic (
    input [1:0] op,
    input [31:0] A, B,
    output [31:0] Y
    );
        
endmodule
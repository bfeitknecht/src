module HalfAdder(input a, input b, output c, output y);

and CARRY(a, b, c);
xor SUM(a, b, y);

endmodule
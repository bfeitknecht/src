module OneTwoDec (
    input s,
    output [1:0] o
);
    // wire ns;
    // not NOTSEL(s, ns);
    // assign o[0] = ns;
    // assign o[1] = s;
endmodule